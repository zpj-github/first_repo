`timescale 1ns/1ps

module add
(


)
ti
od

endmodule
